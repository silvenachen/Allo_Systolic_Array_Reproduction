
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "df_fifo_interface.svh"
`include "df_fifo_monitor.svh"
`include "df_process_interface.svh"
`include "df_process_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "df_loop_interface.svh"
`include "df_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);

    df_fifo_intf fifo_intf_1(clock,reset);
    assign fifo_intf_1.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.indvars_iv26_c_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.indvars_iv26_c_U.if_empty_n;
    assign fifo_intf_1.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.indvars_iv26_c_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.indvars_iv26_c_U.if_full_n;
    assign fifo_intf_1.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.indvars_iv26_blk_n);
    assign fifo_intf_1.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.indvars_iv26_c_blk_n);
    assign fifo_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_1;
    csv_file_dump cstatus_csv_dumper_1;
    df_fifo_monitor fifo_monitor_1;
    df_fifo_intf fifo_intf_2(clock,reset);
    assign fifo_intf_2.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_7_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_7_U.if_empty_n;
    assign fifo_intf_2.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_7_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_7_U.if_full_n;
    assign fifo_intf_2.fifo_rd_block = 0;
    assign fifo_intf_2.fifo_wr_block = 0;
    assign fifo_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_2;
    csv_file_dump cstatus_csv_dumper_2;
    df_fifo_monitor fifo_monitor_2;
    df_fifo_intf fifo_intf_3(clock,reset);
    assign fifo_intf_3.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_6_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_6_U.if_empty_n;
    assign fifo_intf_3.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_6_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_6_U.if_full_n;
    assign fifo_intf_3.fifo_rd_block = 0;
    assign fifo_intf_3.fifo_wr_block = 0;
    assign fifo_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_3;
    csv_file_dump cstatus_csv_dumper_3;
    df_fifo_monitor fifo_monitor_3;
    df_fifo_intf fifo_intf_4(clock,reset);
    assign fifo_intf_4.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_5_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_5_U.if_empty_n;
    assign fifo_intf_4.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_5_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_5_U.if_full_n;
    assign fifo_intf_4.fifo_rd_block = 0;
    assign fifo_intf_4.fifo_wr_block = 0;
    assign fifo_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_4;
    csv_file_dump cstatus_csv_dumper_4;
    df_fifo_monitor fifo_monitor_4;
    df_fifo_intf fifo_intf_5(clock,reset);
    assign fifo_intf_5.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_4_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_4_U.if_empty_n;
    assign fifo_intf_5.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_4_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_4_U.if_full_n;
    assign fifo_intf_5.fifo_rd_block = 0;
    assign fifo_intf_5.fifo_wr_block = 0;
    assign fifo_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_5;
    csv_file_dump cstatus_csv_dumper_5;
    df_fifo_monitor fifo_monitor_5;
    df_fifo_intf fifo_intf_6(clock,reset);
    assign fifo_intf_6.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_3_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_3_U.if_empty_n;
    assign fifo_intf_6.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_3_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_3_U.if_full_n;
    assign fifo_intf_6.fifo_rd_block = 0;
    assign fifo_intf_6.fifo_wr_block = 0;
    assign fifo_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_6;
    csv_file_dump cstatus_csv_dumper_6;
    df_fifo_monitor fifo_monitor_6;
    df_fifo_intf fifo_intf_7(clock,reset);
    assign fifo_intf_7.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_2_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_2_U.if_empty_n;
    assign fifo_intf_7.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_2_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_2_U.if_full_n;
    assign fifo_intf_7.fifo_rd_block = 0;
    assign fifo_intf_7.fifo_wr_block = 0;
    assign fifo_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_7;
    csv_file_dump cstatus_csv_dumper_7;
    df_fifo_monitor fifo_monitor_7;
    df_fifo_intf fifo_intf_8(clock,reset);
    assign fifo_intf_8.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_1_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_1_U.if_empty_n;
    assign fifo_intf_8.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_1_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_1_U.if_full_n;
    assign fifo_intf_8.fifo_rd_block = 0;
    assign fifo_intf_8.fifo_wr_block = 0;
    assign fifo_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_8;
    csv_file_dump cstatus_csv_dumper_8;
    df_fifo_monitor fifo_monitor_8;
    df_fifo_intf fifo_intf_9(clock,reset);
    assign fifo_intf_9.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_U.if_empty_n;
    assign fifo_intf_9.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_C_0_U.if_full_n;
    assign fifo_intf_9.fifo_rd_block = 0;
    assign fifo_intf_9.fifo_wr_block = 0;
    assign fifo_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_9;
    csv_file_dump cstatus_csv_dumper_9;
    df_fifo_monitor fifo_monitor_9;
    df_fifo_intf fifo_intf_10(clock,reset);
    assign fifo_intf_10.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_U.if_empty_n;
    assign fifo_intf_10.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_U.if_full_n;
    assign fifo_intf_10.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.A_fifo_0_blk_n);
    assign fifo_intf_10.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.A_fifo_blk_n);
    assign fifo_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_10;
    csv_file_dump cstatus_csv_dumper_10;
    df_fifo_monitor fifo_monitor_10;
    df_fifo_intf fifo_intf_11(clock,reset);
    assign fifo_intf_11.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_U.if_empty_n;
    assign fifo_intf_11.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_U.if_full_n;
    assign fifo_intf_11.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.B_fifo_0_0_blk_n);
    assign fifo_intf_11.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_blk_n);
    assign fifo_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_11;
    csv_file_dump cstatus_csv_dumper_11;
    df_fifo_monitor fifo_monitor_11;
    df_fifo_intf fifo_intf_12(clock,reset);
    assign fifo_intf_12.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_2_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_2_U.if_empty_n;
    assign fifo_intf_12.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_2_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_2_U.if_full_n;
    assign fifo_intf_12.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.B_fifo_1_0_blk_n);
    assign fifo_intf_12.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_2_blk_n);
    assign fifo_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_12;
    csv_file_dump cstatus_csv_dumper_12;
    df_fifo_monitor fifo_monitor_12;
    df_fifo_intf fifo_intf_13(clock,reset);
    assign fifo_intf_13.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_4_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_4_U.if_empty_n;
    assign fifo_intf_13.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_4_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_4_U.if_full_n;
    assign fifo_intf_13.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.B_fifo_2_0_blk_n);
    assign fifo_intf_13.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_4_blk_n);
    assign fifo_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_13;
    csv_file_dump cstatus_csv_dumper_13;
    df_fifo_monitor fifo_monitor_13;
    df_fifo_intf fifo_intf_14(clock,reset);
    assign fifo_intf_14.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_6_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_6_U.if_empty_n;
    assign fifo_intf_14.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_6_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_6_U.if_full_n;
    assign fifo_intf_14.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.B_fifo_3_0_blk_n);
    assign fifo_intf_14.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_6_blk_n);
    assign fifo_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_14;
    csv_file_dump cstatus_csv_dumper_14;
    df_fifo_monitor fifo_monitor_14;
    df_fifo_intf fifo_intf_15(clock,reset);
    assign fifo_intf_15.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_8_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_8_U.if_empty_n;
    assign fifo_intf_15.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_8_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_8_U.if_full_n;
    assign fifo_intf_15.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.B_fifo_4_0_blk_n);
    assign fifo_intf_15.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_8_blk_n);
    assign fifo_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_15;
    csv_file_dump cstatus_csv_dumper_15;
    df_fifo_monitor fifo_monitor_15;
    df_fifo_intf fifo_intf_16(clock,reset);
    assign fifo_intf_16.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_10_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_10_U.if_empty_n;
    assign fifo_intf_16.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_10_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_10_U.if_full_n;
    assign fifo_intf_16.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.B_fifo_5_0_blk_n);
    assign fifo_intf_16.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_10_blk_n);
    assign fifo_intf_16.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_16;
    csv_file_dump cstatus_csv_dumper_16;
    df_fifo_monitor fifo_monitor_16;
    df_fifo_intf fifo_intf_17(clock,reset);
    assign fifo_intf_17.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_12_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_12_U.if_empty_n;
    assign fifo_intf_17.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_12_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_12_U.if_full_n;
    assign fifo_intf_17.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.B_fifo_6_0_blk_n);
    assign fifo_intf_17.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_12_blk_n);
    assign fifo_intf_17.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_17;
    csv_file_dump cstatus_csv_dumper_17;
    df_fifo_monitor fifo_monitor_17;
    df_fifo_intf fifo_intf_18(clock,reset);
    assign fifo_intf_18.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_14_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_14_U.if_empty_n;
    assign fifo_intf_18.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_14_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_14_U.if_full_n;
    assign fifo_intf_18.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.B_fifo_7_0_blk_n);
    assign fifo_intf_18.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_14_blk_n);
    assign fifo_intf_18.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_18;
    csv_file_dump cstatus_csv_dumper_18;
    df_fifo_monitor fifo_monitor_18;
    df_fifo_intf fifo_intf_19(clock,reset);
    assign fifo_intf_19.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_1_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_1_U.if_empty_n;
    assign fifo_intf_19.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_1_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_1_U.if_full_n;
    assign fifo_intf_19.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.A_fifo_1_blk_n);
    assign fifo_intf_19.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.A_fifo_1_blk_n);
    assign fifo_intf_19.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_19;
    csv_file_dump cstatus_csv_dumper_19;
    df_fifo_monitor fifo_monitor_19;
    df_fifo_intf fifo_intf_20(clock,reset);
    assign fifo_intf_20.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_1_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_1_U.if_empty_n;
    assign fifo_intf_20.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_1_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_1_U.if_full_n;
    assign fifo_intf_20.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_1_blk_n);
    assign fifo_intf_20.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.B_fifo_0_1_blk_n);
    assign fifo_intf_20.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_20;
    csv_file_dump cstatus_csv_dumper_20;
    df_fifo_monitor fifo_monitor_20;
    df_fifo_intf fifo_intf_21(clock,reset);
    assign fifo_intf_21.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_2_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_2_U.if_empty_n;
    assign fifo_intf_21.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_2_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_2_U.if_full_n;
    assign fifo_intf_21.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.A_fifo_2_blk_n);
    assign fifo_intf_21.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.A_fifo_2_blk_n);
    assign fifo_intf_21.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_21;
    csv_file_dump cstatus_csv_dumper_21;
    df_fifo_monitor fifo_monitor_21;
    df_fifo_intf fifo_intf_22(clock,reset);
    assign fifo_intf_22.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_3_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_3_U.if_empty_n;
    assign fifo_intf_22.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_3_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_3_U.if_full_n;
    assign fifo_intf_22.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_3_blk_n);
    assign fifo_intf_22.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.B_fifo_1_1_blk_n);
    assign fifo_intf_22.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_22;
    csv_file_dump cstatus_csv_dumper_22;
    df_fifo_monitor fifo_monitor_22;
    df_fifo_intf fifo_intf_23(clock,reset);
    assign fifo_intf_23.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_3_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_3_U.if_empty_n;
    assign fifo_intf_23.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_3_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_3_U.if_full_n;
    assign fifo_intf_23.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.A_fifo_3_blk_n);
    assign fifo_intf_23.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.A_fifo_3_blk_n);
    assign fifo_intf_23.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_23;
    csv_file_dump cstatus_csv_dumper_23;
    df_fifo_monitor fifo_monitor_23;
    df_fifo_intf fifo_intf_24(clock,reset);
    assign fifo_intf_24.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_5_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_5_U.if_empty_n;
    assign fifo_intf_24.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_5_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_5_U.if_full_n;
    assign fifo_intf_24.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_5_blk_n);
    assign fifo_intf_24.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.B_fifo_2_1_blk_n);
    assign fifo_intf_24.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_24;
    csv_file_dump cstatus_csv_dumper_24;
    df_fifo_monitor fifo_monitor_24;
    df_fifo_intf fifo_intf_25(clock,reset);
    assign fifo_intf_25.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_4_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_4_U.if_empty_n;
    assign fifo_intf_25.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_4_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_4_U.if_full_n;
    assign fifo_intf_25.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.A_fifo_4_blk_n);
    assign fifo_intf_25.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.A_fifo_4_blk_n);
    assign fifo_intf_25.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_25;
    csv_file_dump cstatus_csv_dumper_25;
    df_fifo_monitor fifo_monitor_25;
    df_fifo_intf fifo_intf_26(clock,reset);
    assign fifo_intf_26.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_7_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_7_U.if_empty_n;
    assign fifo_intf_26.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_7_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_7_U.if_full_n;
    assign fifo_intf_26.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_7_blk_n);
    assign fifo_intf_26.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.B_fifo_3_1_blk_n);
    assign fifo_intf_26.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_26;
    csv_file_dump cstatus_csv_dumper_26;
    df_fifo_monitor fifo_monitor_26;
    df_fifo_intf fifo_intf_27(clock,reset);
    assign fifo_intf_27.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_5_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_5_U.if_empty_n;
    assign fifo_intf_27.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_5_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_5_U.if_full_n;
    assign fifo_intf_27.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.A_fifo_5_blk_n);
    assign fifo_intf_27.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.A_fifo_5_blk_n);
    assign fifo_intf_27.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_27;
    csv_file_dump cstatus_csv_dumper_27;
    df_fifo_monitor fifo_monitor_27;
    df_fifo_intf fifo_intf_28(clock,reset);
    assign fifo_intf_28.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_9_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_9_U.if_empty_n;
    assign fifo_intf_28.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_9_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_9_U.if_full_n;
    assign fifo_intf_28.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_9_blk_n);
    assign fifo_intf_28.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.B_fifo_4_1_blk_n);
    assign fifo_intf_28.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_28;
    csv_file_dump cstatus_csv_dumper_28;
    df_fifo_monitor fifo_monitor_28;
    df_fifo_intf fifo_intf_29(clock,reset);
    assign fifo_intf_29.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_6_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_6_U.if_empty_n;
    assign fifo_intf_29.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_6_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_6_U.if_full_n;
    assign fifo_intf_29.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.A_fifo_6_blk_n);
    assign fifo_intf_29.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.A_fifo_6_blk_n);
    assign fifo_intf_29.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_29;
    csv_file_dump cstatus_csv_dumper_29;
    df_fifo_monitor fifo_monitor_29;
    df_fifo_intf fifo_intf_30(clock,reset);
    assign fifo_intf_30.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_11_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_11_U.if_empty_n;
    assign fifo_intf_30.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_11_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_11_U.if_full_n;
    assign fifo_intf_30.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_11_blk_n);
    assign fifo_intf_30.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.B_fifo_5_1_blk_n);
    assign fifo_intf_30.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_30;
    csv_file_dump cstatus_csv_dumper_30;
    df_fifo_monitor fifo_monitor_30;
    df_fifo_intf fifo_intf_31(clock,reset);
    assign fifo_intf_31.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_7_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_7_U.if_empty_n;
    assign fifo_intf_31.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_7_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_7_U.if_full_n;
    assign fifo_intf_31.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.A_fifo_7_blk_n);
    assign fifo_intf_31.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.A_fifo_7_blk_n);
    assign fifo_intf_31.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_31;
    csv_file_dump cstatus_csv_dumper_31;
    df_fifo_monitor fifo_monitor_31;
    df_fifo_intf fifo_intf_32(clock,reset);
    assign fifo_intf_32.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_13_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_13_U.if_empty_n;
    assign fifo_intf_32.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_13_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_13_U.if_full_n;
    assign fifo_intf_32.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_13_blk_n);
    assign fifo_intf_32.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.B_fifo_6_1_blk_n);
    assign fifo_intf_32.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_32;
    csv_file_dump cstatus_csv_dumper_32;
    df_fifo_monitor fifo_monitor_32;
    df_fifo_intf fifo_intf_33(clock,reset);
    assign fifo_intf_33.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_8_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_8_U.if_empty_n;
    assign fifo_intf_33.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_8_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.A_fifo_8_U.if_full_n;
    assign fifo_intf_33.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.A_fifo_8_blk_n);
    assign fifo_intf_33.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.A_fifo_8_blk_n);
    assign fifo_intf_33.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_33;
    csv_file_dump cstatus_csv_dumper_33;
    df_fifo_monitor fifo_monitor_33;
    df_fifo_intf fifo_intf_34(clock,reset);
    assign fifo_intf_34.rd_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_15_U.if_read & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_15_U.if_empty_n;
    assign fifo_intf_34.wr_en = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_15_U.if_write & AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.B_fifo_15_U.if_full_n;
    assign fifo_intf_34.fifo_rd_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_15_blk_n);
    assign fifo_intf_34.fifo_wr_block = ~(AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.B_fifo_7_1_blk_n);
    assign fifo_intf_34.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump fifo_csv_dumper_34;
    csv_file_dump cstatus_csv_dumper_34;
    df_fifo_monitor fifo_monitor_34;

logic region_0_idle;
logic [31:0] region_0_start_cnt;
logic [31:0] region_0_done_cnt;
assign region_0_idle = (region_0_start_cnt == region_0_done_cnt) && AESL_inst_systolic_modulate.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_start_cnt <= 32'h0;
    else if (AESL_inst_systolic_modulate.ap_start == 1'b1 && AESL_inst_systolic_modulate.ap_ready == 1'b1)
        region_0_start_cnt <= region_0_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_0_done_cnt <= 32'h0;
    else if (AESL_inst_systolic_modulate.ap_done == 1'b1)
        region_0_done_cnt <= region_0_done_cnt + 32'h1;
    else;
end

logic region_1_idle;
logic [31:0] region_1_start_cnt;
logic [31:0] region_1_done_cnt;
assign region_1_idle = (region_1_start_cnt == region_1_done_cnt) && AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_start_cnt <= 32'h0;
    else if (AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_start == 1'b1 && AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_ready == 1'b1)
        region_1_start_cnt <= region_1_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_1_done_cnt <= 32'h0;
    else if (AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_done == 1'b1 && AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_continue == 1'b1)
        region_1_done_cnt <= region_1_done_cnt + 32'h1;
    else;
end

logic region_2_idle;
logic [31:0] region_2_start_cnt;
logic [31:0] region_2_done_cnt;
assign region_2_idle = (region_2_start_cnt == region_2_done_cnt) && AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_start == 1'b0 ;
always @(posedge clock) begin
    if (reset == 1'b1)
        region_2_start_cnt <= 32'h0;
    else if (AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_start == 1'b1 && AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_ready == 1'b1)
        region_2_start_cnt <= region_2_start_cnt + 32'h1;
    else;
end
always @(posedge clock) begin
    if (reset == 1'b1)
        region_2_done_cnt <= 32'h0;
    else if (AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_done == 1'b1 && AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_continue == 1'b1)
        region_2_done_cnt <= region_2_done_cnt + 32'h1;
    else;
end


    df_process_intf process_intf_1(clock,reset);
    assign process_intf_1.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_start;
    assign process_intf_1.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_ready;
    assign process_intf_1.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_done;
    assign process_intf_1.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_continue;
    assign process_intf_1.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_start;
    assign process_intf_1.pin_stall = 1'b0;
    assign process_intf_1.pout_stall = 1'b0;
    assign process_intf_1.cin_stall = 1'b0;
    assign process_intf_1.cout_stall = 1'b0;
    assign process_intf_1.region_idle = region_0_idle;
    assign process_intf_1.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_1;
    csv_file_dump pstatus_csv_dumper_1;
    df_process_monitor process_monitor_1;
    df_process_intf process_intf_2(clock,reset);
    assign process_intf_2.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.ap_start;
    assign process_intf_2.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.ap_ready;
    assign process_intf_2.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.ap_done;
    assign process_intf_2.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.ap_continue;
    assign process_intf_2.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.ap_start;
    assign process_intf_2.pin_stall = 1'b0;
    assign process_intf_2.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.indvars_iv26_c_blk_n;
    assign process_intf_2.cin_stall = 1'b0;
    assign process_intf_2.cout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_A_0_U.i_full_n;
    assign process_intf_2.region_idle = region_1_idle;
    assign process_intf_2.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_2;
    csv_file_dump pstatus_csv_dumper_2;
    df_process_monitor process_monitor_2;
    df_process_intf process_intf_3(clock,reset);
    assign process_intf_3.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_start;
    assign process_intf_3.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_ready;
    assign process_intf_3.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_done;
    assign process_intf_3.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_continue;
    assign process_intf_3.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_start;
    assign process_intf_3.pin_stall = 1'b0;
    assign process_intf_3.pout_stall = 1'b0;
    assign process_intf_3.cin_stall = 1'b0;
    assign process_intf_3.cout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_1_49_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_2_50_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_3_51_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_3_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_2_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_1_U.i_full_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_4_U.i_full_n;
    assign process_intf_3.region_idle = region_1_idle;
    assign process_intf_3.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_3;
    csv_file_dump pstatus_csv_dumper_3;
    df_process_monitor process_monitor_3;
    df_process_intf process_intf_4(clock,reset);
    assign process_intf_4.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_start;
    assign process_intf_4.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_ready;
    assign process_intf_4.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_done;
    assign process_intf_4.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_continue;
    assign process_intf_4.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.ap_start;
    assign process_intf_4.pin_stall = 1'b0;
    assign process_intf_4.pout_stall = 1'b0;
    assign process_intf_4.cin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_A_0_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_4_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_1_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_2_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_3_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_3_51_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_2_50_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_1_49_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_U.t_empty_n;
    assign process_intf_4.cout_stall = 1'b0;
    assign process_intf_4.region_idle = region_1_idle;
    assign process_intf_4.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_4;
    csv_file_dump pstatus_csv_dumper_4;
    df_process_monitor process_monitor_4;
    df_process_intf process_intf_5(clock,reset);
    assign process_intf_5.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_start;
    assign process_intf_5.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_ready;
    assign process_intf_5.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_done;
    assign process_intf_5.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_continue;
    assign process_intf_5.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.real_start;
    assign process_intf_5.pin_stall = 1'b0;
    assign process_intf_5.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.A_fifo_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_2_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_4_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_6_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_8_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_10_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_12_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.B_fifo_14_blk_n;
    assign process_intf_5.cin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_A_0_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_4_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_1_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_2_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_3_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_3_51_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_2_50_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_1_49_U.t_empty_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.local_B_U.t_empty_n;
    assign process_intf_5.cout_stall = 1'b0;
    assign process_intf_5.region_idle = region_2_idle;
    assign process_intf_5.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_5;
    csv_file_dump pstatus_csv_dumper_5;
    df_process_monitor process_monitor_5;
    df_process_intf process_intf_6(clock,reset);
    assign process_intf_6.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_start;
    assign process_intf_6.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_ready;
    assign process_intf_6.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_done;
    assign process_intf_6.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_continue;
    assign process_intf_6.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.real_start;
    assign process_intf_6.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.A_fifo_0_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.B_fifo_0_0_blk_n;
    assign process_intf_6.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.A_fifo_1_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.B_fifo_0_1_blk_n;
    assign process_intf_6.cin_stall = 1'b0;
    assign process_intf_6.cout_stall = 1'b0;
    assign process_intf_6.region_idle = region_2_idle;
    assign process_intf_6.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_6;
    csv_file_dump pstatus_csv_dumper_6;
    df_process_monitor process_monitor_6;
    df_process_intf process_intf_7(clock,reset);
    assign process_intf_7.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_start;
    assign process_intf_7.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_ready;
    assign process_intf_7.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_done;
    assign process_intf_7.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_continue;
    assign process_intf_7.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_start;
    assign process_intf_7.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.A_fifo_1_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.B_fifo_1_0_blk_n;
    assign process_intf_7.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.A_fifo_2_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.B_fifo_1_1_blk_n;
    assign process_intf_7.cin_stall = 1'b0;
    assign process_intf_7.cout_stall = 1'b0;
    assign process_intf_7.region_idle = region_2_idle;
    assign process_intf_7.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_7;
    csv_file_dump pstatus_csv_dumper_7;
    df_process_monitor process_monitor_7;
    df_process_intf process_intf_8(clock,reset);
    assign process_intf_8.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_start;
    assign process_intf_8.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_ready;
    assign process_intf_8.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_done;
    assign process_intf_8.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_continue;
    assign process_intf_8.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_start;
    assign process_intf_8.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.A_fifo_2_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.B_fifo_2_0_blk_n;
    assign process_intf_8.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.A_fifo_3_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.B_fifo_2_1_blk_n;
    assign process_intf_8.cin_stall = 1'b0;
    assign process_intf_8.cout_stall = 1'b0;
    assign process_intf_8.region_idle = region_2_idle;
    assign process_intf_8.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_8;
    csv_file_dump pstatus_csv_dumper_8;
    df_process_monitor process_monitor_8;
    df_process_intf process_intf_9(clock,reset);
    assign process_intf_9.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_start;
    assign process_intf_9.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_ready;
    assign process_intf_9.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_done;
    assign process_intf_9.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_continue;
    assign process_intf_9.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_start;
    assign process_intf_9.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.A_fifo_3_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.B_fifo_3_0_blk_n;
    assign process_intf_9.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.A_fifo_4_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.B_fifo_3_1_blk_n;
    assign process_intf_9.cin_stall = 1'b0;
    assign process_intf_9.cout_stall = 1'b0;
    assign process_intf_9.region_idle = region_2_idle;
    assign process_intf_9.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_9;
    csv_file_dump pstatus_csv_dumper_9;
    df_process_monitor process_monitor_9;
    df_process_intf process_intf_10(clock,reset);
    assign process_intf_10.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_start;
    assign process_intf_10.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_ready;
    assign process_intf_10.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_done;
    assign process_intf_10.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_continue;
    assign process_intf_10.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_start;
    assign process_intf_10.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.A_fifo_4_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.B_fifo_4_0_blk_n;
    assign process_intf_10.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.A_fifo_5_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.B_fifo_4_1_blk_n;
    assign process_intf_10.cin_stall = 1'b0;
    assign process_intf_10.cout_stall = 1'b0;
    assign process_intf_10.region_idle = region_2_idle;
    assign process_intf_10.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_10;
    csv_file_dump pstatus_csv_dumper_10;
    df_process_monitor process_monitor_10;
    df_process_intf process_intf_11(clock,reset);
    assign process_intf_11.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_start;
    assign process_intf_11.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_ready;
    assign process_intf_11.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_done;
    assign process_intf_11.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_continue;
    assign process_intf_11.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_start;
    assign process_intf_11.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.A_fifo_5_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.B_fifo_5_0_blk_n;
    assign process_intf_11.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.A_fifo_6_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.B_fifo_5_1_blk_n;
    assign process_intf_11.cin_stall = 1'b0;
    assign process_intf_11.cout_stall = 1'b0;
    assign process_intf_11.region_idle = region_2_idle;
    assign process_intf_11.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_11;
    csv_file_dump pstatus_csv_dumper_11;
    df_process_monitor process_monitor_11;
    df_process_intf process_intf_12(clock,reset);
    assign process_intf_12.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_start;
    assign process_intf_12.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_ready;
    assign process_intf_12.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_done;
    assign process_intf_12.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_continue;
    assign process_intf_12.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_start;
    assign process_intf_12.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.A_fifo_6_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.B_fifo_6_0_blk_n;
    assign process_intf_12.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.A_fifo_7_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.B_fifo_6_1_blk_n;
    assign process_intf_12.cin_stall = 1'b0;
    assign process_intf_12.cout_stall = 1'b0;
    assign process_intf_12.region_idle = region_2_idle;
    assign process_intf_12.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_12;
    csv_file_dump pstatus_csv_dumper_12;
    df_process_monitor process_monitor_12;
    df_process_intf process_intf_13(clock,reset);
    assign process_intf_13.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_start;
    assign process_intf_13.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_ready;
    assign process_intf_13.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_done;
    assign process_intf_13.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_continue;
    assign process_intf_13.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_start;
    assign process_intf_13.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.A_fifo_7_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.B_fifo_7_0_blk_n;
    assign process_intf_13.pout_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.A_fifo_8_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.B_fifo_7_1_blk_n;
    assign process_intf_13.cin_stall = 1'b0;
    assign process_intf_13.cout_stall = 1'b0;
    assign process_intf_13.region_idle = region_2_idle;
    assign process_intf_13.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_13;
    csv_file_dump pstatus_csv_dumper_13;
    df_process_monitor process_monitor_13;
    df_process_intf process_intf_14(clock,reset);
    assign process_intf_14.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_start;
    assign process_intf_14.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_ready;
    assign process_intf_14.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_done;
    assign process_intf_14.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_continue;
    assign process_intf_14.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_start;
    assign process_intf_14.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.A_fifo_8_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_1_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_3_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_5_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_7_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_9_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_11_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_13_blk_n | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.B_fifo_15_blk_n;
    assign process_intf_14.pout_stall = 1'b0;
    assign process_intf_14.cin_stall = 1'b0;
    assign process_intf_14.cout_stall = 1'b0;
    assign process_intf_14.region_idle = region_2_idle;
    assign process_intf_14.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_14;
    csv_file_dump pstatus_csv_dumper_14;
    df_process_monitor process_monitor_14;
    df_process_intf process_intf_15(clock,reset);
    assign process_intf_15.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.ap_start;
    assign process_intf_15.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.ap_ready;
    assign process_intf_15.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.ap_done;
    assign process_intf_15.ap_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.ap_continue;
    assign process_intf_15.real_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.ap_start;
    assign process_intf_15.pin_stall = 1'b0 | ~AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.indvars_iv26_blk_n;
    assign process_intf_15.pout_stall = 1'b0;
    assign process_intf_15.cin_stall = 1'b0;
    assign process_intf_15.cout_stall = 1'b0;
    assign process_intf_15.region_idle = region_1_idle;
    assign process_intf_15.finish = finish | deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock;
    csv_file_dump pstall_csv_dumper_15;
    csv_file_dump pstatus_csv_dumper_15;
    df_process_monitor process_monitor_15;

    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_systolic_modulate.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_systolic_modulate.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_systolic_modulate.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;

    pp_loop_intf #(4) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_1.post_states_valid = 1'b1;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_1.quit_at_end = 1'b1;
    assign pp_loop_intf_1.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_0_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(4) pp_loop_monitor_1;
    pp_loop_intf #(4) pp_loop_intf_2(clock,reset);
    assign pp_loop_intf_2.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_2.pre_states_valid = 1'b1;
    assign pp_loop_intf_2.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_2.post_states_valid = 1'b1;
    assign pp_loop_intf_2.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_2.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_2.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_2.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_2.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_2.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_2.quit_at_end = 1'b1;
    assign pp_loop_intf_2.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_1_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_2.finish = finish;
    csv_file_dump pp_loop_csv_dumper_2;
    pp_loop_monitor #(4) pp_loop_monitor_2;
    pp_loop_intf #(4) pp_loop_intf_3(clock,reset);
    assign pp_loop_intf_3.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_3.pre_states_valid = 1'b1;
    assign pp_loop_intf_3.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_3.post_states_valid = 1'b1;
    assign pp_loop_intf_3.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_3.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_3.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_3.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_3.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_3.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_3.quit_at_end = 1'b1;
    assign pp_loop_intf_3.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_2_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_3.finish = finish;
    csv_file_dump pp_loop_csv_dumper_3;
    pp_loop_monitor #(4) pp_loop_monitor_3;
    pp_loop_intf #(4) pp_loop_intf_4(clock,reset);
    assign pp_loop_intf_4.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_4.pre_states_valid = 1'b1;
    assign pp_loop_intf_4.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_4.post_states_valid = 1'b1;
    assign pp_loop_intf_4.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_4.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_4.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_4.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_4.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_4.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_4.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_4.quit_at_end = 1'b1;
    assign pp_loop_intf_4.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_3_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_4.finish = finish;
    csv_file_dump pp_loop_csv_dumper_4;
    pp_loop_monitor #(4) pp_loop_monitor_4;
    pp_loop_intf #(4) pp_loop_intf_5(clock,reset);
    assign pp_loop_intf_5.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_5.pre_states_valid = 1'b1;
    assign pp_loop_intf_5.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_5.post_states_valid = 1'b1;
    assign pp_loop_intf_5.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_5.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_5.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_5.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_5.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_5.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_5.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_5.quit_at_end = 1'b1;
    assign pp_loop_intf_5.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_4_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_5.finish = finish;
    csv_file_dump pp_loop_csv_dumper_5;
    pp_loop_monitor #(4) pp_loop_monitor_5;
    pp_loop_intf #(4) pp_loop_intf_6(clock,reset);
    assign pp_loop_intf_6.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_6.pre_states_valid = 1'b1;
    assign pp_loop_intf_6.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_6.post_states_valid = 1'b1;
    assign pp_loop_intf_6.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_6.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_6.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_6.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_6.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_6.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_6.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_6.quit_at_end = 1'b1;
    assign pp_loop_intf_6.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_5_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_6.finish = finish;
    csv_file_dump pp_loop_csv_dumper_6;
    pp_loop_monitor #(4) pp_loop_monitor_6;
    pp_loop_intf #(4) pp_loop_intf_7(clock,reset);
    assign pp_loop_intf_7.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_7.pre_states_valid = 1'b1;
    assign pp_loop_intf_7.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_7.post_states_valid = 1'b1;
    assign pp_loop_intf_7.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_7.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_7.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_7.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_7.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_7.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_7.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_7.quit_at_end = 1'b1;
    assign pp_loop_intf_7.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_6_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_7.finish = finish;
    csv_file_dump pp_loop_csv_dumper_7;
    pp_loop_monitor #(4) pp_loop_monitor_7;
    pp_loop_intf #(4) pp_loop_intf_8(clock,reset);
    assign pp_loop_intf_8.pre_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_ST_fsm_state1;
    assign pp_loop_intf_8.pre_states_valid = 1'b1;
    assign pp_loop_intf_8.post_loop_state0 = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_ST_fsm_state8;
    assign pp_loop_intf_8.post_states_valid = 1'b1;
    assign pp_loop_intf_8.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_8.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_8.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_8.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_8.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_enable_reg_pp0_iter2;
    assign pp_loop_intf_8.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_block_pp0_stage1_subdone;
    assign pp_loop_intf_8.loop_quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_ST_fsm_pp0_stage1;
    assign pp_loop_intf_8.quit_at_end = 1'b1;
    assign pp_loop_intf_8.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.PE_kernel_modulate_7_0_1_U0.ap_CS_fsm;
    assign pp_loop_intf_8.finish = finish;
    csv_file_dump pp_loop_csv_dumper_8;
    pp_loop_monitor #(4) pp_loop_monitor_8;
    df_loop_intf df_loop_intf_1(clock,reset);
    assign df_loop_intf_1.body_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_start;
    assign df_loop_intf_1.body_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_ready;
    assign df_loop_intf_1.body_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_done;
    assign df_loop_intf_1.body_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.ap_continue;
    assign df_loop_intf_1.loop_start = AESL_inst_systolic_modulate.ap_start;
    assign df_loop_intf_1.loop_ready = AESL_inst_systolic_modulate.ap_ready;
    assign df_loop_intf_1.loop_done = AESL_inst_systolic_modulate.ap_done;
    assign df_loop_intf_1.loop_continue = 1'b1;
    csv_file_dump df_loop_csv_dumper_1;
    df_loop_monitor df_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.loop_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_load_A_tile_ak_proc_Pipeline_l_load_A_tile_ak_fu_50.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;
    upc_loop_intf#(1) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.quit_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.loop_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_done;
    assign upc_loop_intf_2.loop_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_load_B_tile_bk_proc_U0.ap_continue;
    assign upc_loop_intf_2.quit_at_end = 1'b1;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(1) upc_loop_monitor_2;
    upc_loop_intf#(1) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.quit_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_3.loop_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_done;
    assign upc_loop_intf_3.loop_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_load_k8_proc21_U0.ap_continue;
    assign upc_loop_intf_3.quit_at_end = 1'b1;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(1) upc_loop_monitor_3;
    upc_loop_intf#(1) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.quit_enable = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.loop_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_done;
    assign upc_loop_intf_4.loop_continue = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.systolic_tile_modulate_U0.systolic_tile_modulate_Loop_l_data_drain_k9_proc22_U0.ap_continue;
    assign upc_loop_intf_4.quit_at_end = 1'b1;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(1) upc_loop_monitor_4;
    upc_loop_intf#(1) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ST_fsm_state1;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ST_fsm_state1;
    assign upc_loop_intf_5.quit_state = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ST_fsm_state1;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_5.quit_block = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ST_fsm_state1_blk;
    assign upc_loop_intf_5.iter_start_enable = 1'b1;
    assign upc_loop_intf_5.iter_end_enable = 1'b1;
    assign upc_loop_intf_5.quit_enable = 1'b1;
    assign upc_loop_intf_5.loop_start = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_systolic_modulate.dataflow_in_loop_l_ni_1_U0.dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_U0.grp_dataflow_in_loop_l_ni_1_Loop_l_store_C_tile_sj_proc_Pipeline_l_store_C_tile_sj_fu_104.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b1;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(1) upc_loop_monitor_5;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;

    fifo_csv_dumper_1 = new("./depth1.csv");
    cstatus_csv_dumper_1 = new("./chan_status1.csv");
    fifo_monitor_1 = new(fifo_csv_dumper_1,fifo_intf_1,cstatus_csv_dumper_1);
    fifo_csv_dumper_2 = new("./depth2.csv");
    cstatus_csv_dumper_2 = new("./chan_status2.csv");
    fifo_monitor_2 = new(fifo_csv_dumper_2,fifo_intf_2,cstatus_csv_dumper_2);
    fifo_csv_dumper_3 = new("./depth3.csv");
    cstatus_csv_dumper_3 = new("./chan_status3.csv");
    fifo_monitor_3 = new(fifo_csv_dumper_3,fifo_intf_3,cstatus_csv_dumper_3);
    fifo_csv_dumper_4 = new("./depth4.csv");
    cstatus_csv_dumper_4 = new("./chan_status4.csv");
    fifo_monitor_4 = new(fifo_csv_dumper_4,fifo_intf_4,cstatus_csv_dumper_4);
    fifo_csv_dumper_5 = new("./depth5.csv");
    cstatus_csv_dumper_5 = new("./chan_status5.csv");
    fifo_monitor_5 = new(fifo_csv_dumper_5,fifo_intf_5,cstatus_csv_dumper_5);
    fifo_csv_dumper_6 = new("./depth6.csv");
    cstatus_csv_dumper_6 = new("./chan_status6.csv");
    fifo_monitor_6 = new(fifo_csv_dumper_6,fifo_intf_6,cstatus_csv_dumper_6);
    fifo_csv_dumper_7 = new("./depth7.csv");
    cstatus_csv_dumper_7 = new("./chan_status7.csv");
    fifo_monitor_7 = new(fifo_csv_dumper_7,fifo_intf_7,cstatus_csv_dumper_7);
    fifo_csv_dumper_8 = new("./depth8.csv");
    cstatus_csv_dumper_8 = new("./chan_status8.csv");
    fifo_monitor_8 = new(fifo_csv_dumper_8,fifo_intf_8,cstatus_csv_dumper_8);
    fifo_csv_dumper_9 = new("./depth9.csv");
    cstatus_csv_dumper_9 = new("./chan_status9.csv");
    fifo_monitor_9 = new(fifo_csv_dumper_9,fifo_intf_9,cstatus_csv_dumper_9);
    fifo_csv_dumper_10 = new("./depth10.csv");
    cstatus_csv_dumper_10 = new("./chan_status10.csv");
    fifo_monitor_10 = new(fifo_csv_dumper_10,fifo_intf_10,cstatus_csv_dumper_10);
    fifo_csv_dumper_11 = new("./depth11.csv");
    cstatus_csv_dumper_11 = new("./chan_status11.csv");
    fifo_monitor_11 = new(fifo_csv_dumper_11,fifo_intf_11,cstatus_csv_dumper_11);
    fifo_csv_dumper_12 = new("./depth12.csv");
    cstatus_csv_dumper_12 = new("./chan_status12.csv");
    fifo_monitor_12 = new(fifo_csv_dumper_12,fifo_intf_12,cstatus_csv_dumper_12);
    fifo_csv_dumper_13 = new("./depth13.csv");
    cstatus_csv_dumper_13 = new("./chan_status13.csv");
    fifo_monitor_13 = new(fifo_csv_dumper_13,fifo_intf_13,cstatus_csv_dumper_13);
    fifo_csv_dumper_14 = new("./depth14.csv");
    cstatus_csv_dumper_14 = new("./chan_status14.csv");
    fifo_monitor_14 = new(fifo_csv_dumper_14,fifo_intf_14,cstatus_csv_dumper_14);
    fifo_csv_dumper_15 = new("./depth15.csv");
    cstatus_csv_dumper_15 = new("./chan_status15.csv");
    fifo_monitor_15 = new(fifo_csv_dumper_15,fifo_intf_15,cstatus_csv_dumper_15);
    fifo_csv_dumper_16 = new("./depth16.csv");
    cstatus_csv_dumper_16 = new("./chan_status16.csv");
    fifo_monitor_16 = new(fifo_csv_dumper_16,fifo_intf_16,cstatus_csv_dumper_16);
    fifo_csv_dumper_17 = new("./depth17.csv");
    cstatus_csv_dumper_17 = new("./chan_status17.csv");
    fifo_monitor_17 = new(fifo_csv_dumper_17,fifo_intf_17,cstatus_csv_dumper_17);
    fifo_csv_dumper_18 = new("./depth18.csv");
    cstatus_csv_dumper_18 = new("./chan_status18.csv");
    fifo_monitor_18 = new(fifo_csv_dumper_18,fifo_intf_18,cstatus_csv_dumper_18);
    fifo_csv_dumper_19 = new("./depth19.csv");
    cstatus_csv_dumper_19 = new("./chan_status19.csv");
    fifo_monitor_19 = new(fifo_csv_dumper_19,fifo_intf_19,cstatus_csv_dumper_19);
    fifo_csv_dumper_20 = new("./depth20.csv");
    cstatus_csv_dumper_20 = new("./chan_status20.csv");
    fifo_monitor_20 = new(fifo_csv_dumper_20,fifo_intf_20,cstatus_csv_dumper_20);
    fifo_csv_dumper_21 = new("./depth21.csv");
    cstatus_csv_dumper_21 = new("./chan_status21.csv");
    fifo_monitor_21 = new(fifo_csv_dumper_21,fifo_intf_21,cstatus_csv_dumper_21);
    fifo_csv_dumper_22 = new("./depth22.csv");
    cstatus_csv_dumper_22 = new("./chan_status22.csv");
    fifo_monitor_22 = new(fifo_csv_dumper_22,fifo_intf_22,cstatus_csv_dumper_22);
    fifo_csv_dumper_23 = new("./depth23.csv");
    cstatus_csv_dumper_23 = new("./chan_status23.csv");
    fifo_monitor_23 = new(fifo_csv_dumper_23,fifo_intf_23,cstatus_csv_dumper_23);
    fifo_csv_dumper_24 = new("./depth24.csv");
    cstatus_csv_dumper_24 = new("./chan_status24.csv");
    fifo_monitor_24 = new(fifo_csv_dumper_24,fifo_intf_24,cstatus_csv_dumper_24);
    fifo_csv_dumper_25 = new("./depth25.csv");
    cstatus_csv_dumper_25 = new("./chan_status25.csv");
    fifo_monitor_25 = new(fifo_csv_dumper_25,fifo_intf_25,cstatus_csv_dumper_25);
    fifo_csv_dumper_26 = new("./depth26.csv");
    cstatus_csv_dumper_26 = new("./chan_status26.csv");
    fifo_monitor_26 = new(fifo_csv_dumper_26,fifo_intf_26,cstatus_csv_dumper_26);
    fifo_csv_dumper_27 = new("./depth27.csv");
    cstatus_csv_dumper_27 = new("./chan_status27.csv");
    fifo_monitor_27 = new(fifo_csv_dumper_27,fifo_intf_27,cstatus_csv_dumper_27);
    fifo_csv_dumper_28 = new("./depth28.csv");
    cstatus_csv_dumper_28 = new("./chan_status28.csv");
    fifo_monitor_28 = new(fifo_csv_dumper_28,fifo_intf_28,cstatus_csv_dumper_28);
    fifo_csv_dumper_29 = new("./depth29.csv");
    cstatus_csv_dumper_29 = new("./chan_status29.csv");
    fifo_monitor_29 = new(fifo_csv_dumper_29,fifo_intf_29,cstatus_csv_dumper_29);
    fifo_csv_dumper_30 = new("./depth30.csv");
    cstatus_csv_dumper_30 = new("./chan_status30.csv");
    fifo_monitor_30 = new(fifo_csv_dumper_30,fifo_intf_30,cstatus_csv_dumper_30);
    fifo_csv_dumper_31 = new("./depth31.csv");
    cstatus_csv_dumper_31 = new("./chan_status31.csv");
    fifo_monitor_31 = new(fifo_csv_dumper_31,fifo_intf_31,cstatus_csv_dumper_31);
    fifo_csv_dumper_32 = new("./depth32.csv");
    cstatus_csv_dumper_32 = new("./chan_status32.csv");
    fifo_monitor_32 = new(fifo_csv_dumper_32,fifo_intf_32,cstatus_csv_dumper_32);
    fifo_csv_dumper_33 = new("./depth33.csv");
    cstatus_csv_dumper_33 = new("./chan_status33.csv");
    fifo_monitor_33 = new(fifo_csv_dumper_33,fifo_intf_33,cstatus_csv_dumper_33);
    fifo_csv_dumper_34 = new("./depth34.csv");
    cstatus_csv_dumper_34 = new("./chan_status34.csv");
    fifo_monitor_34 = new(fifo_csv_dumper_34,fifo_intf_34,cstatus_csv_dumper_34);

    pstall_csv_dumper_1 = new("./stalling1.csv");
    pstatus_csv_dumper_1 = new("./status1.csv");
    process_monitor_1 = new(pstall_csv_dumper_1,process_intf_1,pstatus_csv_dumper_1);
    pstall_csv_dumper_2 = new("./stalling2.csv");
    pstatus_csv_dumper_2 = new("./status2.csv");
    process_monitor_2 = new(pstall_csv_dumper_2,process_intf_2,pstatus_csv_dumper_2);
    pstall_csv_dumper_3 = new("./stalling3.csv");
    pstatus_csv_dumper_3 = new("./status3.csv");
    process_monitor_3 = new(pstall_csv_dumper_3,process_intf_3,pstatus_csv_dumper_3);
    pstall_csv_dumper_4 = new("./stalling4.csv");
    pstatus_csv_dumper_4 = new("./status4.csv");
    process_monitor_4 = new(pstall_csv_dumper_4,process_intf_4,pstatus_csv_dumper_4);
    pstall_csv_dumper_5 = new("./stalling5.csv");
    pstatus_csv_dumper_5 = new("./status5.csv");
    process_monitor_5 = new(pstall_csv_dumper_5,process_intf_5,pstatus_csv_dumper_5);
    pstall_csv_dumper_6 = new("./stalling6.csv");
    pstatus_csv_dumper_6 = new("./status6.csv");
    process_monitor_6 = new(pstall_csv_dumper_6,process_intf_6,pstatus_csv_dumper_6);
    pstall_csv_dumper_7 = new("./stalling7.csv");
    pstatus_csv_dumper_7 = new("./status7.csv");
    process_monitor_7 = new(pstall_csv_dumper_7,process_intf_7,pstatus_csv_dumper_7);
    pstall_csv_dumper_8 = new("./stalling8.csv");
    pstatus_csv_dumper_8 = new("./status8.csv");
    process_monitor_8 = new(pstall_csv_dumper_8,process_intf_8,pstatus_csv_dumper_8);
    pstall_csv_dumper_9 = new("./stalling9.csv");
    pstatus_csv_dumper_9 = new("./status9.csv");
    process_monitor_9 = new(pstall_csv_dumper_9,process_intf_9,pstatus_csv_dumper_9);
    pstall_csv_dumper_10 = new("./stalling10.csv");
    pstatus_csv_dumper_10 = new("./status10.csv");
    process_monitor_10 = new(pstall_csv_dumper_10,process_intf_10,pstatus_csv_dumper_10);
    pstall_csv_dumper_11 = new("./stalling11.csv");
    pstatus_csv_dumper_11 = new("./status11.csv");
    process_monitor_11 = new(pstall_csv_dumper_11,process_intf_11,pstatus_csv_dumper_11);
    pstall_csv_dumper_12 = new("./stalling12.csv");
    pstatus_csv_dumper_12 = new("./status12.csv");
    process_monitor_12 = new(pstall_csv_dumper_12,process_intf_12,pstatus_csv_dumper_12);
    pstall_csv_dumper_13 = new("./stalling13.csv");
    pstatus_csv_dumper_13 = new("./status13.csv");
    process_monitor_13 = new(pstall_csv_dumper_13,process_intf_13,pstatus_csv_dumper_13);
    pstall_csv_dumper_14 = new("./stalling14.csv");
    pstatus_csv_dumper_14 = new("./status14.csv");
    process_monitor_14 = new(pstall_csv_dumper_14,process_intf_14,pstatus_csv_dumper_14);
    pstall_csv_dumper_15 = new("./stalling15.csv");
    pstatus_csv_dumper_15 = new("./status15.csv");
    process_monitor_15 = new(pstall_csv_dumper_15,process_intf_15,pstatus_csv_dumper_15);

    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);
    pp_loop_csv_dumper_2 = new("./pp_loop_status2.csv");
    pp_loop_monitor_2 = new(pp_loop_intf_2,pp_loop_csv_dumper_2);
    pp_loop_csv_dumper_3 = new("./pp_loop_status3.csv");
    pp_loop_monitor_3 = new(pp_loop_intf_3,pp_loop_csv_dumper_3);
    pp_loop_csv_dumper_4 = new("./pp_loop_status4.csv");
    pp_loop_monitor_4 = new(pp_loop_intf_4,pp_loop_csv_dumper_4);
    pp_loop_csv_dumper_5 = new("./pp_loop_status5.csv");
    pp_loop_monitor_5 = new(pp_loop_intf_5,pp_loop_csv_dumper_5);
    pp_loop_csv_dumper_6 = new("./pp_loop_status6.csv");
    pp_loop_monitor_6 = new(pp_loop_intf_6,pp_loop_csv_dumper_6);
    pp_loop_csv_dumper_7 = new("./pp_loop_status7.csv");
    pp_loop_monitor_7 = new(pp_loop_intf_7,pp_loop_csv_dumper_7);
    pp_loop_csv_dumper_8 = new("./pp_loop_status8.csv");
    pp_loop_monitor_8 = new(pp_loop_intf_8,pp_loop_csv_dumper_8);
    df_loop_csv_dumper_1 = new("./df_loop_status1.csv");
    df_loop_monitor_1 = new(df_loop_intf_1,df_loop_csv_dumper_1);



    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);

    sample_manager_inst.add_one_monitor(fifo_monitor_1);
    sample_manager_inst.add_one_monitor(fifo_monitor_2);
    sample_manager_inst.add_one_monitor(fifo_monitor_3);
    sample_manager_inst.add_one_monitor(fifo_monitor_4);
    sample_manager_inst.add_one_monitor(fifo_monitor_5);
    sample_manager_inst.add_one_monitor(fifo_monitor_6);
    sample_manager_inst.add_one_monitor(fifo_monitor_7);
    sample_manager_inst.add_one_monitor(fifo_monitor_8);
    sample_manager_inst.add_one_monitor(fifo_monitor_9);
    sample_manager_inst.add_one_monitor(fifo_monitor_10);
    sample_manager_inst.add_one_monitor(fifo_monitor_11);
    sample_manager_inst.add_one_monitor(fifo_monitor_12);
    sample_manager_inst.add_one_monitor(fifo_monitor_13);
    sample_manager_inst.add_one_monitor(fifo_monitor_14);
    sample_manager_inst.add_one_monitor(fifo_monitor_15);
    sample_manager_inst.add_one_monitor(fifo_monitor_16);
    sample_manager_inst.add_one_monitor(fifo_monitor_17);
    sample_manager_inst.add_one_monitor(fifo_monitor_18);
    sample_manager_inst.add_one_monitor(fifo_monitor_19);
    sample_manager_inst.add_one_monitor(fifo_monitor_20);
    sample_manager_inst.add_one_monitor(fifo_monitor_21);
    sample_manager_inst.add_one_monitor(fifo_monitor_22);
    sample_manager_inst.add_one_monitor(fifo_monitor_23);
    sample_manager_inst.add_one_monitor(fifo_monitor_24);
    sample_manager_inst.add_one_monitor(fifo_monitor_25);
    sample_manager_inst.add_one_monitor(fifo_monitor_26);
    sample_manager_inst.add_one_monitor(fifo_monitor_27);
    sample_manager_inst.add_one_monitor(fifo_monitor_28);
    sample_manager_inst.add_one_monitor(fifo_monitor_29);
    sample_manager_inst.add_one_monitor(fifo_monitor_30);
    sample_manager_inst.add_one_monitor(fifo_monitor_31);
    sample_manager_inst.add_one_monitor(fifo_monitor_32);
    sample_manager_inst.add_one_monitor(fifo_monitor_33);
    sample_manager_inst.add_one_monitor(fifo_monitor_34);
    sample_manager_inst.add_one_monitor(process_monitor_1);
    sample_manager_inst.add_one_monitor(process_monitor_2);
    sample_manager_inst.add_one_monitor(process_monitor_3);
    sample_manager_inst.add_one_monitor(process_monitor_4);
    sample_manager_inst.add_one_monitor(process_monitor_5);
    sample_manager_inst.add_one_monitor(process_monitor_6);
    sample_manager_inst.add_one_monitor(process_monitor_7);
    sample_manager_inst.add_one_monitor(process_monitor_8);
    sample_manager_inst.add_one_monitor(process_monitor_9);
    sample_manager_inst.add_one_monitor(process_monitor_10);
    sample_manager_inst.add_one_monitor(process_monitor_11);
    sample_manager_inst.add_one_monitor(process_monitor_12);
    sample_manager_inst.add_one_monitor(process_monitor_13);
    sample_manager_inst.add_one_monitor(process_monitor_14);
    sample_manager_inst.add_one_monitor(process_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_2);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_3);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_4);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_5);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_6);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_7);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_8);
    sample_manager_inst.add_one_monitor(df_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1 || deadlock_detector.AESL_deadlock_report_unit_inst.find_df_deadlock == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
